// Copyright (C) 2022  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 21.1.1 Build 850 06/23/2022 SJ Lite Edition"
// CREATED		"Tue Aug 15 19:23:26 2023"

module CMP2(
	A,
	B,
	G,
	E,
	L
);


input wire	[1:0] A;
input wire	[1:0] B;
output wire	G;
output wire	E;
output wire	L;

wire	E_ALTERA_SYNTHESIZED0;
wire	E_ALTERA_SYNTHESIZED1;
wire	G_ALTERA_SYNTHESIZED0;
wire	G_ALTERA_SYNTHESIZED1;
wire	L_ALTERA_SYNTHESIZED0;
wire	L_ALTERA_SYNTHESIZED1;
wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;




assign	G = SYNTHESIZED_WIRE_0 | G_ALTERA_SYNTHESIZED1;


CMP1	b2v_inst1(
	.A(A[1]),
	.B(B[1]),
	.G(G_ALTERA_SYNTHESIZED1),
	.E(E_ALTERA_SYNTHESIZED1),
	.L(L_ALTERA_SYNTHESIZED1));


CMP1	b2v_inst2(
	.A(A[0]),
	.B(B[0]),
	.G(G_ALTERA_SYNTHESIZED0),
	.E(E_ALTERA_SYNTHESIZED0),
	.L(L_ALTERA_SYNTHESIZED0));

assign	SYNTHESIZED_WIRE_0 = E_ALTERA_SYNTHESIZED1 & G_ALTERA_SYNTHESIZED0;

assign	L = SYNTHESIZED_WIRE_1 | L_ALTERA_SYNTHESIZED1;

assign	SYNTHESIZED_WIRE_1 = E_ALTERA_SYNTHESIZED1 & L_ALTERA_SYNTHESIZED0;

assign	E = E_ALTERA_SYNTHESIZED1 & E_ALTERA_SYNTHESIZED0;


endmodule
